LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY circuito2 IS
	PORT (
		A2, A1, A0 								: IN STD_LOGIC;
		S0, S1, S2, S3, S4, S5, S6, S7 	: OUT STD_LOGIC
	);
END circuito2;

ARCHITECTURE behavior OF circuito2 IS
BEGIN
	S0 <= '1' WHEN (NOT A2 AND NOT A1 AND NOT A0) = '1' ELSE '0';
	S1 <= '1' WHEN (NOT A2 AND NOT A1 AND A0) = '1' ELSE '0';
	S2 <= '1' WHEN (NOT A2 AND A1 AND NOT A0) = '1' ELSE '0';
	S3 <= '1' WHEN (NOT A2 AND A1 AND A0) = '1' ELSE '0';
	S4 <= '1' WHEN (A2 AND NOT A1 AND NOT A0) = '1' ELSE '0';
	S5 <= '1' WHEN (A2 AND NOT A1 AND A0) = '1' ELSE '0';
	S6 <= '1' WHEN (A2 AND A1 AND NOT A0) = '1' ELSE '0';
	S7 <= '1' WHEN (A2 AND A1 AND A0) = '1' ELSE '0';
END behavior;