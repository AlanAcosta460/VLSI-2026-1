LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY circuito3 IS
	PORT (
		A2, A1, A0 								: IN STD_LOGIC;
		S0, S1, S2, S3, S4, S5, S6, S7 	: OUT STD_LOGIC
	);
END circuito3;

ARCHITECTURE behavior OF circuito3 IS
BEGIN
	WITH (NOT A2 AND NOT A1 AND NOT A0) SELECT
		S0 <= '1' WHEN '1',
				'0' WHEN OTHERS;
	
	WITH (NOT A2 AND NOT A1 AND A0) SELECT
		S1 <= '1' WHEN '1',
				'0' WHEN OTHERS;
	
	WITH (NOT A2 AND A1 AND NOT A0) SELECT
		S2 <= '1' WHEN '1',
				'0' WHEN OTHERS;
		
	WITH (NOT A2 AND A1 AND A0) SELECT
		S3 <= '1' WHEN '1',
				'0' WHEN OTHERS;
		
	WITH (A2 AND NOT A1 AND NOT A0) SELECT
		S4 <= '1' WHEN '1',
				'0' WHEN OTHERS;
		
	WITH (A2 AND NOT A1 AND A0) SELECT
		S5 <= '1' WHEN '1',
				'0' WHEN OTHERS;
		
	WITH (A2 AND A1 AND NOT A0) SELECT
		S6 <= '1' WHEN '1',
				'0' WHEN OTHERS;
		
	WITH (A2 AND A1 AND A0) SELECT
		S7 <= '1' WHEN '1',
				'0' WHEN OTHERS;
END behavior;