LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY circuito1 IS
    PORT (
        D3, D2, D1, D0             : IN STD_LOGIC;
        Sa, Sb, Sc, Sd, Se, Sf, Sg : OUT STD_LOGIC
    );
END circuito1;

ARCHITECTURE behavior OF circuito1 IS
BEGIN
    Sa <= (NOT D3 AND D1) OR
          (NOT D3 AND NOT D2 AND NOT D0) OR
          (NOT D3 AND D2 AND D0) OR
          (D3 AND NOT D2 AND NOT D1);
            
    Sb <= (NOT D3 AND NOT D2) OR
          (NOT D2 AND NOT D1) OR
          (NOT D3 AND NOT D1 AND NOT D0) OR
          (NOT D3 AND D1 AND D0);
            
    Sc <= (NOT D2 AND NOT D1) OR
          (NOT D3 AND D0) OR
          (NOT D3 AND D2);
            
    Sd <= (NOT D2 AND NOT D1 AND NOT D0) OR
          (NOT D3 AND NOT D2 AND D1) OR
          (NOT D3 AND D1 AND NOT D0) OR
          (NOT D3 AND D2 AND NOT D1 AND D0);
            
    Se <= (NOT D2 AND NOT D1 AND NOT D0) OR
          (NOT D3 AND D1 AND NOT D0);
            
    Sf <= (NOT D2 AND NOT D1 AND NOT D0) OR
          (NOT D3 AND D2 AND NOT D0) OR
          (NOT D3 AND D2 AND NOT D1) OR
          (D3 AND NOT D2 AND NOT D1);
            
    Sg <= (NOT D3 AND NOT D2 AND D1) OR
          (NOT D3 AND D2 AND NOT D0) OR
          (NOT D3 AND D2 AND NOT D1) OR
          (D3 AND NOT D2 AND NOT D1);
END behavior;
