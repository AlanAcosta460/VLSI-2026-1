LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY and_1 IS PORT(
	I1, I2	: IN STD_LOGIC;
	O1			: OUT STD_LOGIC
);
END and_1;

ARCHITECTURE dataflow OF and_1 IS
BEGIN
	O1 <= I1 AND I2;
end dataflow;


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY or_1 IS PORT(
	I1, I2	: IN STD_LOGIC;
	O1			: OUT STD_LOGIC
);
END or_1;

ARCHITECTURE dataflow OF or_1 IS
BEGIN
	O1 <= I1 OR I2;
end dataflow;


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY xor_1 IS PORT(
	I1, I2	: IN STD_LOGIC;
	O1			: OUT STD_LOGIC
);
END xor_1;

ARCHITECTURE dataflow OF xor_1 IS
BEGIN
	O1 <= I1 XOR I2;
end dataflow;


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY nand_1 IS PORT(
	I1, I2	: IN STD_LOGIC;
	O1			: OUT STD_LOGIC
);
END nand_1;

ARCHITECTURE dataflow OF nand_1 IS
BEGIN
	O1 <= NOT(I1 AND I2);
end dataflow;


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY xnor_1 IS PORT(
	I1, I2	: IN STD_LOGIC;
	O1			: OUT STD_LOGIC
);
END xnor_1;

ARCHITECTURE dataflow OF xnor_1 IS
BEGIN
	O1 <= NOT(I1 XOR I2);
end dataflow;


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY circuito2 IS PORT(
	A, B, C	: IN STD_LOGIC;
	S1, S2	: OUT STD_LOGIC
);
END circuito2;

ARCHITECTURE structural OF circuito2 IS
	SIGNAL Y1, Y2, Y3, Y4 : STD_LOGIC;
	
	COMPONENT and_1 IS PORT(
		I1, I2	: IN STD_LOGIC;
		O1			: OUT STD_LOGIC
	);
	END COMPONENT;
	
	COMPONENT or_1 IS PORT(
		I1, I2	: IN STD_LOGIC;
		O1			: OUT STD_LOGIC
	);
	END COMPONENT;
	
	COMPONENT xor_1 IS PORT(
		I1, I2	: IN STD_LOGIC;
		O1			: OUT STD_LOGIC
	);
	END COMPONENT;
	
	COMPONENT nand_1 IS PORT(
		I1, I2	: IN STD_LOGIC;
		O1			: OUT STD_LOGIC
	);
	END COMPONENT;
	
	COMPONENT xnor_1 IS PORT(
		I1, I2	: IN STD_LOGIC;
		O1			: OUT STD_LOGIC
	);
	END COMPONENT;
BEGIN
	C1: xnor_1 PORT MAP(I1 => A, I2 => B, O1 => Y1);
	C2: xor_1 PORT MAP(I1 => Y1, I2 => C, O1 => S1);
	
	C3: nand_1 PORT MAP(I1 => A, I2 => B, O1 => Y2);
	C4: or_1 PORT MAP(I1 => A, I2 => B, O1 => Y3);
	C5: and_1 PORT MAP(I1 => Y3, I2 => C, O1 => Y4);
	C6: or_1 PORT MAP(I1 => Y2, I2 => Y4, O1 => S2);
END structural;
