LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY circuito7 IS PORT (
    A, B, C             : IN STD_LOGIC;
    S1A, S2A, S1B, S2B  : OUT STD_LOGIC
);
END circuito7;

ARCHITECTURE arc OF circuito7 IS
	SIGNAL Y1, Y2, Y3, Y4 : STD_LOGIC;
BEGIN
	S1A <= (A XNOR B) XOR C;
	S2A <= (A NAND B) OR ((A OR B) AND C);

	proceso: PROCESS (A, B, C)
	BEGIN
		Y1 <= A XNOR B;
		S1B <= Y1 XOR C;
		
		Y2 <= A NAND B;
		Y3 <= A OR B;
		Y4 <= Y3 AND C;
		S2B <= Y2 OR Y4;
	END PROCESS proceso;
END arc;
