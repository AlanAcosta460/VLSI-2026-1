LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY circuito1 IS
	PORT (
		A2, A1, A0 								: IN STD_LOGIC;
		S0, S1, S2, S3, S4, S5, S6, S7 	: OUT STD_LOGIC
	);
END circuito1;

ARCHITECTURE behavior OF circuito1 IS
BEGIN
	S0 <= NOT A2 AND NOT A1 AND NOT A0;
	S1 <= NOT A2 AND NOT A1 AND A0;
	S2 <= NOT A2 AND A1 AND NOT A0;
	S3 <= NOT A2 AND A1 AND A0;
	S4 <= A2 AND NOT A1 AND NOT A0;
	S5 <= A2 AND NOT A1 AND A0;
	S6 <= A2 AND A1 AND NOT A0;
	S7 <= A2 AND A1 AND A0;
END behavior;