LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY and_1 IS PORT(
	I1, I2	: IN STD_LOGIC;
	O1			: OUT STD_LOGIC
);
END and_1;

ARCHITECTURE dataflow OF and_1 IS
BEGIN
	O1 <= I1 AND I2;
end dataflow;


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY or_1 IS PORT(
	I1, I2	: IN STD_LOGIC;
	O1			: OUT STD_LOGIC
);
END or_1;

ARCHITECTURE dataflow OF or_1 IS
BEGIN
	O1 <= I1 OR I2;
end dataflow;


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY nor_1 IS PORT(
	I1, I2	: IN STD_LOGIC;
	O1			: OUT STD_LOGIC
);
END nor_1;

ARCHITECTURE dataflow OF nor_1 IS
BEGIN
	O1 <= NOT(I1 OR I2);
end dataflow;


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY xnor_1 IS PORT(
	I1, I2	: IN STD_LOGIC;
	O1			: OUT STD_LOGIC
);
END xnor_1;

ARCHITECTURE dataflow OF xnor_1 IS
BEGIN
	O1 <= NOT(I1 XOR I2);
end dataflow;


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY circuito1 IS PORT(
	A, B, C	: IN STD_LOGIC;
	F, E		: OUT STD_LOGIC
);
END circuito1;

ARCHITECTURE structural OF circuito1 IS
	SIGNAL Y1, Y2, Y3, Y4 : STD_LOGIC;
	
	COMPONENT and_1 IS PORT(
		I1, I2	: IN STD_LOGIC;
		O1			: OUT STD_LOGIC
	);
	END COMPONENT;
	
	COMPONENT or_1 IS PORT(
		I1, I2	: IN STD_LOGIC;
		O1			: OUT STD_LOGIC
	);
	END COMPONENT;
	
	COMPONENT nor_1 IS PORT(
		I1, I2	: IN STD_LOGIC;
		O1			: OUT STD_LOGIC
	);
	END COMPONENT;
	
	COMPONENT xnor_1 IS PORT(
		I1, I2	: IN STD_LOGIC;
		O1			: OUT STD_LOGIC
	);
	END COMPONENT;
BEGIN
	C1: and_1 PORT MAP(I1 => A, I2 => B, O1 => Y1);
	C2: and_1 PORT MAP(I1 => B, I2 => C, O1 => Y2);
	C3: xnor_1 PORT MAP(I1 => Y1, I2 => Y2, O1 => Y3);
	C4: or_1 PORT MAP(I1 => A, I2 => Y3, O1 => F);
	
	C5: nor_1 PORT MAP(I1 => A, I2 => Y2, O1 => Y4);
	C6: or_1 PORT MAP(I1 => Y4, I2 => C, O1 => E);
END structural;
